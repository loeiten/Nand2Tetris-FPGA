`default_nettype none
module Hack2(
    input clk_in,				// external clock 100 MHz
    input [7:0] but,			// buttons	(0 if pressed, 1 if released)
    output [7:0] led,			// LEDs 	(0 off, 1 on)
    input rx,					// rx line of UART
    output tx					// tx line of UART
  );





endmodule
