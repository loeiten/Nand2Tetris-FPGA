/**
 * 16-bit Not:
 * for i=0..15: out[i] = not in[i]
 */
`default_nettype none

module Not16(
    input [15:0] in,
    output [15:0] out
  );



endmodule
