/**
 * 16-bit bitwise And:
 * for i = 0..15: out[i] = (a[i] and b[i])
 */

`default_nettype none
module And16(
    input wire [15:0] a,
    input wire [15:0] b,
    output wire [15:0] out
  );

  // your implementation comes here:



endmodule
