`default_nettype none
module Hack1(
    input clk_in,				// external clock 100 MHz
    input [1:0] but,			// buttons	(0 if pressed, 1 if released)
	output [1:0] led			// leds 	(0 off, 1 on)
);




endmodule
