/**
* Timer
*
* real time module increments out[16] by one every 0.0001 seconds.
* doesn't care about overflow.
*/

`default_nettype none
module Timer(
    input wire clk,
    output wire [15:0] out
  );




endmodule
